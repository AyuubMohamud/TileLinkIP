module i2cphy();
endmodule
