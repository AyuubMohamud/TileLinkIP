module openPolarisI2C (
    
);
    
endmodule
