module polaris_dma
#(
    parameter NoC = 2 //! Number of channels to generate
)
(
    
);
    
endmodule
