module DMACore (
    
);
    
endmodule
