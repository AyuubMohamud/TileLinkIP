//! TileLink many masters to 1 slave (Non-blocking)