module spiphy (
    
);
    
endmodule